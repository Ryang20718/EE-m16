//--------------------------------------------------------------------
//		Timescale
//		Means that if you do #1 in the initial block of your
//		testbench, time is advanced by 1ns instead of 1ps
//--------------------------------------------------------------------
`timescale 1ns / 1ps

//--------------------------------------------------------------------
//		Design Assign #2, Testbench.
//--------------------------------------------------------------------
//
// This is a model of the motor for you to test the motor drive signal. It includes a count to see if the position is correct
//
module motor(count, err, motor_drv, drv_clk, reset);
   output [7:0]    count;
   output 	err;
   input [3:0] 	motor_drv;
   input 	drv_clk, reset;

   reg signed [7:0] count;
   reg 		err;
   reg [3:0] 	prev_motor_drv;
   
   always @(motor_drv or reset) begin
      if (reset) begin
	 count = 0;
	 prev_motor_drv=4'b0000;
      end
      else begin
	 case (motor_drv)
	   4'b0000: begin
	      // $display("No Motor Drive: drv=%b prev_drv=%b", motor_drv, prev_motor_drv);
	   end
	   4'b0001: begin
	      err = 0;
	      if (prev_motor_drv == 4'b0010)
		count = count-1;
	      else if (prev_motor_drv == 4'b1000)
		count = count+1;
	      else if (prev_motor_drv == 4'b0001)
		;
	      // $display("No Motor Change: drv=%b prev_drv=%b", motor_drv, prev_motor_drv);		
	      else if (prev_motor_drv == 4'b0000)
		;
	      // $display("From Reset: drv=%b prev_drv=%b", motor_drv, prev_motor_drv);		
	      else begin
		 // $display("ERR: drv=%b prev_drv=%b", motor_drv, prev_motor_drv);
		 err = 1;
	      end
	      prev_motor_drv=4'b0001;
	   end
	   4'b0011: begin
	      if ((prev_motor_drv!==4'b0001) || (prev_motor_drv!==4'b0010)) begin
		 // $display("ERR: drv=%b prev_drv=%b", motor_drv, prev_motor_drv);
		 err = 1;
	      end
	   end
	   4'b0010: begin
	      err = 0;
	      if (prev_motor_drv == 4'b0100)
		count = count-1;
	      else if (prev_motor_drv == 4'b0001)
		count = count+1;
	      else if (prev_motor_drv == 4'b0010)
		;
  	      // $display("No Motor Change: drv=%b prev_drv=%b", motor_drv, prev_motor_drv);		
	      else begin
		 // $display("ERR: drv=%b prev_drv=%b", motor_drv, prev_motor_drv);
		 err = 1;
	      end
	      prev_motor_drv=4'b0010;
	   end
	   4'b0110: begin
      	      if ((prev_motor_drv!==4'b0100) || (prev_motor_drv!==4'b0010)) begin
		 // $display("ERR: drv=%b prev_drv=%b", motor_drv, prev_motor_drv);
		 err = 1;
	      end
	   end
	   4'b0100: begin
	      err = 0;
	      if (prev_motor_drv == 4'b1000)
		count = count-1;
	      else if (prev_motor_drv == 4'b0010)
		count = count+1;
	      else if (prev_motor_drv == 4'b0100)
		;
	      // $display("No Motor Change: drv=%b prev_drv=%b", motor_drv, prev_motor_drv);		
	      else begin
		 // $display("ERR: drv=%b prev_drv=%b", motor_drv, prev_motor_drv);
		 err = 1;
	      end
	      prev_motor_drv=4'b0100;
	   end
	   4'b1100: begin
      	      if ((prev_motor_drv!==4'b1000) || (prev_motor_drv!==4'b0001)) begin
		 // $display("ERR: drv=%b prev_drv=%b", motor_drv, prev_motor_drv);
		 err = 1;
	      end
	   end
	   4'b1000: begin
	      err = 0;
	      if (prev_motor_drv == 4'b0001)
		count = count-1;
	      else if (prev_motor_drv == 4'b0100)
		count = count+1;
	      else if (prev_motor_drv == 4'b1000)
		;
	      // $display("No Change: drv=%b prev_drv=%b", motor_drv, prev_motor_drv);		
	      else begin
		 // $display("ERR: drv=%b prev_drv=%b", motor_drv, prev_motor_drv);
		 err = 1;
	      end
	      prev_motor_drv=4'b1000;
	   end
	   4'b1001: begin
      	      if ((prev_motor_drv!==4'b1000) || (prev_motor_drv!==4'b0001)) begin
		 // $display("ERR: drv=%b prev_drv=%b", motor_drv, prev_motor_drv);
		 err = 1;
	      end
	   end
	   default: begin
	      // $display("ERR: drv=%b prev_drv=%b", motor_drv, prev_motor_drv);
	      err = 1;	      
	   end
	 endcase // case (motor_drv)
      end // else: !if(reset)
   end // always @ (motor_drv or reset)
endmodule // motor

//
// This is the module that generates a clock for you to use in your design
//
module clkgen(clk);
   output clk;

   reg 	  clk;
   
   initial
     clk = 1'b0;
   always
     #100 clk=~clk;
endmodule

module dassign2_tb();
   //----------------------------------------------------------------
   //		Test Bench Signal Declarations
   //----------------------------------------------------------------
   integer i,j,outfile;
   //----------------------------------------------------------------
   //		Instantiate modules Module
   //----------------------------------------------------------------
   clkgen clkgen_1(drv_clk);
   motor motor_1(step_count, step_err, motor_drv, drv_clk, reset);
   
   sbs sbs_tst(diff, bout, in0, in1, bin);
   dassign2_1	dassign2_1(quot, remout, remin, div);
   dassign2_2	dassign2_2(motor_drv, done, forward, reverse, reset, drv_clk);
   //----------------------------------------------------------------
   //		Design Task #1 Signal Declarations
   //----------------------------------------------------------------
   wire    diff, bout;
   reg 	   in0, in1, bin;

   wire    quot;
   wire [7:0] remout;
   reg [7:0]  remin, div;

   reg [8:0]  din0, din1, dout;
   reg [7:0]  tstrem;
   reg 	      tstquot;

   integer    sbs_err, sub_err, scs_err;
   //----------------------------------------------------------------
   //		Design Task #2 Signal Declarations
   //----------------------------------------------------------------
   wire [3:0] motor_drv;
   wire       done, drv_clk;
   reg 	      forward, reverse, reset;

   wire signed [7:0] step_count;
   wire       step_err;
   
   integer    motseq_err, forw_err, rev_err, done_err;
   //----------------------------------------------------------------
   //		Test Stimulus
   //----------------------------------------------------------------
   initial begin
      outfile=$fopen("dassign2.txt");
      if(!outfile) begin
	 $display("FAIL WRITE FILE");
	 $finish;
      end
      $dumpfile("dassign2.vcd");
      $dumpvars(0,dassign2_tb);
      sbs_err = 0;
      sub_err = 0;
      scs_err = 0;
      #1 ;
      din0 = 0;
      din1 = 0;
      #1 ;
      for(i=0;i<8;i=i+1) begin
	 {in0, in1, bin} = i[2:0];
	 #1 ;
	 din0[0] = in0;
	 din1[0] = in1;
	 dout = din0 - din1 - bin;
	 if ((dout[0] !== diff) || (dout[1] !== bout))
	   sbs_err = sbs_err + 1;
	 //      $display(i, in0, in1, bin, diff, bout, din0, din1, dout, dout[0], dout[1]);
      end
      #1 ;
      for(i=0;i<256;i=i+1) begin
	 div[7:0] = i[7:0];
	 #1
	   for(j=0;j<256;j=j+1) begin
	      remin[7:0] = j[7:0];
	      #1 ;
	      dout[8:0] = remin[7:0] - div[7:0];
	      #1 ;
	      if (dout[8] === 1'b1) begin
		 tstquot = 1'b0;
		 tstrem[7:0] = remin[7:0];
	      end
	      else begin
		 tstquot = 1'b1;
		 tstrem[7:0] = dout[7:0];
	      end
	      #1 ;
	      if (dassign2_1.dout !== dout[7:0])
		sub_err = sub_err + 1;
	      if ((tstrem !== remout) || (tstquot !== quot))
		scs_err = scs_err + 1;
	      // $display(i, div, j, remin, "\t", dout[7:0], "\t", dassign2_1.dout, "\t", remout, "\t", tstrem, "\t\t",dout[8], ~quot, sub_err, scs_err);	 
	   end
      end
      $display("SBS ERR: %d", sbs_err);
      $display("Subtractor ERR: %d", sub_err);
      $display("SCS ERR: %d", scs_err);
      #100 ;
      motseq_err = 0;
      forw_err = 0;
      rev_err = 0;
      done_err = 0;
      forward = 0;
      reverse = 0;
      reset = 1;
      #200 ;
      reset = 0;
      for(i=0;i<8;i=i+1) begin
	 forward = 1;
	 #200 ;
	// $display("forw %b\trev %b\tmotor_drv %b\tstep_count %d", forward, reverse, motor_drv, step_count);
         forward = 0;
	 #200 ;
	 // $display("forw %b\trev %b\tmotor_drv %b\tstep_count %d", forward, reverse, motor_drv, step_count);
      end
      if (step_count != 8) begin
	$display("ERR: incorrect position.");
	 forw_err = forw_err+1;
      end
      for(i=0;i<8;i=i+1) begin
	 forward = 1;
	 #200 ;
	 // $display("forw %b\trev %b\tmotor_drv %b\tstep_count %d", forward, reverse, motor_drv, step_count);
      end
      if (step_count != 16) begin
	 $display("ERR: incorrect position.");
	 forw_err = forw_err+1;
      end
      forward = 0;
      #200 ;
      // $display("forw %b\trev %b\tmotor_drv %b\tstep_count %d", forward, reverse, motor_drv, step_count);
      for(i=0;i<32;i=i+1) begin
	 reverse = 1;
	 #200 ;
	 // $display("forw %b\trev %b\tmotor_drv %b\tstep_count %d", forward, reverse, motor_drv, step_count);
      end
      if (step_count != -16) begin
	 $display("ERR: incorrect position.");
	 rev_err = rev_err+1;
      end
      for(i=0;i<16;i=i+1) begin
	 reverse = 1;
	 #200 ;
	 reverse = 0;
	 #200 ;
	 // $display("forw %b\trev %b\tmotor_drv %b\tstep_count %d", forward, reverse, motor_drv, step_count);
      end
      if (step_count != -32) begin
	 $display("ERR: incorrect position.");
	 rev_err = rev_err+1;
      end
      #200;
      #200;
      #200;
      $finish;
   end // initial begin
   always @(posedge drv_clk) begin
      if (done)
	if (step_count %4 == 0)
	  ;
          // $display ("done asserted at step count:", step_count);
	else begin
	   $display ("ERR: done");
	   done_err = done_err + 1;
	end
      if (step_err) begin
	 $display ("ERR: at step count, %d, motor drve %b", step_count, motor_drv);
	 motseq_err = motseq_err + 1;
      end 
   end
endmodule // dassign2_tb


